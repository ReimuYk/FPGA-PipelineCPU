module add4(in,out4);
	input [31:0] in;
	output [31:0] out4;
	
	assign out4 = in+4;
endmodule
