module reg_D(pc4, ins, wpcir, clock, resetn, dpc4, dins);
	input	[31:0]	pc4, ins;
	input				wpcir, clock, resetn;
	output[31:0]	dpc4, dins;
	
	/* need to complete */
endmodule
