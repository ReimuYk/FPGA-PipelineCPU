module reg_W(mwreg, mm2reg, 
malu, mmo, mrn, 
clock, resetn, 
wwreg, wm2reg, wmo, walu, wrn);
	input         mwreg, mm2reg, clock, resetn;
	input  [4:0]  mrn;
	input  [31:0] mmo, malu;
	output        wwreg, wm2reg;
	output [4:0]  wrn;
	output [31:0] wmo, walu;
	
	/* need to complete */
endmodule
